module Ejercicio2(input a,output b);
	assign b=a;
endmodule