module DisplayTest(input a,output b);
	assign b=a;

endmodule